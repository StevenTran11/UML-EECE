-- sim_street_image.vhd
--
-- FPGA Vision Remote Lab http://h-brs.de/fpga-vision-lab
-- (c) Marco Winzker, Hochschule Bonn-Rhein-Sieg, 02.05.2019

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use std.textio.all;
use ieee.std_logic_textio.all;

entity sim_street_image is
end sim_street_image;

architecture sim of sim_street_image is

-- signals of testbench
  signal clk_25    : std_logic := '0';
  signal reset     : std_logic;
  signal vs_out    : std_logic;
  signal hs_out    : std_logic;
  signal de_out    : std_logic;
  signal r_out     : std_logic_vector(7 downto 0);
  signal g_out     : std_logic_vector(7 downto 0);
  signal b_out     : std_logic_vector(7 downto 0);
  
begin

-- clock generation
  clk_25 <= not clk_25 after 20 ns;

-- reset
  reset  <= '1', '0' after 95 ns;
  
  
-- instantiation of design-under-verification
  duv : entity work.street_image
    port map (clk_25        => clk_25,
              reset         => reset,
              vs_out        => vs_out,
              hs_out        => hs_out,
              de_out        => de_out,
              r_out         => r_out,
              g_out         => g_out,
              b_out         => b_out);


-- write output to ppm-file
-- ppm-file can be viewed with IrfanView and probably other image viewers
-- verified with IrfanView version 4.44 - 64 bit
-- EXPERIMENTAL, please give feedback in case of problems

  file_process : process

    file     response_file     : text;
    constant response_filename : string  := "image_out.ppm";
    variable l_o               : line;
    variable response_status   : file_open_status;
    variable x_size            : integer := 640;
    variable y_size            : integer := 480;
    variable x, y              : integer;

  begin

    -- open output file
    file_open(response_status, response_file, response_filename, write_mode);
    write (l_o, string'("P3"));       -- magic number
    writeline(response_file, l_o);        
    write (l_o, string'("# generated by VHDL testbench"));       -- comment
    writeline(response_file, l_o);        
    write (l_o, x_size);
    write (l_o, string'(" "));
    write (l_o, y_size);
    writeline(response_file, l_o);        
    write (l_o, string'("255"));       -- maximum value
    writeline(response_file, l_o);        
        
    -- write pixel to file
    for y in 0 to y_size-1 loop
    wait until rising_edge(de_out); -- begin of line

      for x in 0 to x_size-1 loop
      wait until falling_edge(clk_25); -- middle of clock cycle

        write (l_o, to_integer(unsigned(r_out)));
        write (l_o, string'(" "));
        write (l_o, to_integer(unsigned(g_out)));
        write (l_o, string'(" "));
        write (l_o, to_integer(unsigned(b_out)));
        writeline(response_file, l_o);        
       
        end loop;  -- x
    end loop;  -- y

    wait for 1000 ns;

    file_close(response_file);
    assert false
      report "Simulation completed"
      severity failure;

  end process;


end sim;